module language

pub const grandfathereds = ['i-default', 'i-mingo']
