module tests

struct WithError {
mut:
	error IError
}
