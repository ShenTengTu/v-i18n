module language

pub const extlangs = ['ar-aao', 'ar-abh', 'ar-abv', 'ar-acm', 'ar-acq', 'ar-acw', 'ar-acx', 'ar-acy',
	'ar-adf', 'ar-aeb', 'ar-aec', 'ar-afb', 'ar-ajp', 'ar-apc', 'ar-apd', 'ar-arb', 'ar-arq',
	'ar-ars', 'ar-ary', 'ar-arz', 'ar-auz', 'ar-avl', 'ar-ayh', 'ar-ayl', 'ar-ayn', 'ar-ayp',
	'ar-pga', 'ar-shu', 'ar-ssh', 'kok-gom', 'kok-knn', 'lv-ltg', 'lv-lvs', 'ms-bjn', 'ms-btj',
	'ms-bve', 'ms-bvu', 'ms-coa', 'ms-dup', 'ms-hji', 'ms-jak', 'ms-jax', 'ms-kvb', 'ms-kvr',
	'ms-kxd', 'ms-lce', 'ms-lcf', 'ms-liw', 'ms-max', 'ms-meo', 'ms-mfa', 'ms-mfb', 'ms-min',
	'ms-mqg', 'ms-msi', 'ms-mui', 'ms-orn', 'ms-ors', 'ms-pel', 'ms-pse', 'ms-tmw', 'ms-urk',
	'ms-vkk', 'ms-vkt', 'ms-xmm', 'ms-zlm', 'ms-zmi', 'ms-zsm', 'sgn-ads', 'sgn-aed', 'sgn-aen',
	'sgn-afg', 'sgn-ase', 'sgn-asf', 'sgn-asp', 'sgn-asq', 'sgn-asw', 'sgn-bfi', 'sgn-bfk', 'sgn-bog',
	'sgn-bqn', 'sgn-bqy', 'sgn-bvl', 'sgn-bzs', 'sgn-cds', 'sgn-csc', 'sgn-csd', 'sgn-cse', 'sgn-csf',
	'sgn-csg', 'sgn-csl', 'sgn-csn', 'sgn-csq', 'sgn-csr', 'sgn-csx', 'sgn-doq', 'sgn-dse', 'sgn-dsl',
	'sgn-ecs', 'sgn-ehs', 'sgn-esl', 'sgn-esn', 'sgn-eso', 'sgn-eth', 'sgn-fcs', 'sgn-fse', 'sgn-fsl',
	'sgn-fss', 'sgn-gds', 'sgn-gse', 'sgn-gsg', 'sgn-gsm', 'sgn-gss', 'sgn-gus', 'sgn-hab', 'sgn-haf',
	'sgn-hds', 'sgn-hks', 'sgn-hos', 'sgn-hps', 'sgn-hsh', 'sgn-hsl', 'sgn-icl', 'sgn-iks', 'sgn-ils',
	'sgn-inl', 'sgn-ins', 'sgn-ise', 'sgn-isg', 'sgn-isr', 'sgn-jcs', 'sgn-jhs', 'sgn-jks', 'sgn-jls',
	'sgn-jos', 'sgn-jsl', 'sgn-jus', 'sgn-kgi', 'sgn-kvk', 'sgn-lbs', 'sgn-lls', 'sgn-lsb', 'sgn-lsl',
	'sgn-lsn', 'sgn-lso', 'sgn-lsp', 'sgn-lst', 'sgn-lsv', 'sgn-lsy', 'sgn-lws', 'sgn-mdl', 'sgn-mfs',
	'sgn-mre', 'sgn-msd', 'sgn-msr', 'sgn-mzc', 'sgn-mzg', 'sgn-mzy', 'sgn-nbs', 'sgn-ncs', 'sgn-nsi',
	'sgn-nsl', 'sgn-nsp', 'sgn-nsr', 'sgn-nzs', 'sgn-okl', 'sgn-pgz', 'sgn-pks', 'sgn-prl', 'sgn-prz',
	'sgn-psc', 'sgn-psd', 'sgn-psg', 'sgn-psl', 'sgn-pso', 'sgn-psp', 'sgn-psr', 'sgn-pys', 'sgn-rms',
	'sgn-rsl', 'sgn-rsm', 'sgn-sdl', 'sgn-sfb', 'sgn-sfs', 'sgn-sgg', 'sgn-sgx', 'sgn-slf', 'sgn-sls',
	'sgn-sqk', 'sgn-sqs', 'sgn-sqx', 'sgn-ssp', 'sgn-ssr', 'sgn-svk', 'sgn-swl', 'sgn-syy', 'sgn-szs',
	'sgn-tse', 'sgn-tsm', 'sgn-tsq', 'sgn-tss', 'sgn-tsy', 'sgn-tza', 'sgn-ugn', 'sgn-ugy', 'sgn-ukl',
	'sgn-uks', 'sgn-vgt', 'sgn-vsi', 'sgn-vsl', 'sgn-vsv', 'sgn-wbs', 'sgn-xki', 'sgn-xml', 'sgn-xms',
	'sgn-ygs', 'sgn-yhs', 'sgn-ysl', 'sgn-ysm', 'sgn-zib', 'sgn-zsl', 'sw-swc', 'sw-swh', 'uz-uzn',
	'uz-uzs', 'zh-cdo', 'zh-cjy', 'zh-cmn', 'zh-cnp', 'zh-cpx', 'zh-csp', 'zh-czh', 'zh-czo',
	'zh-gan', 'zh-hak', 'zh-hsn', 'zh-lzh', 'zh-mnp', 'zh-nan', 'zh-wuu', 'zh-yue']
