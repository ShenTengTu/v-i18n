module i18n

const version = '0.0.0-alpha'
