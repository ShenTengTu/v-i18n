module language

pub const redundants = ['az-Arab', 'az-Cyrl', 'az-Latn', 'be-Latn', 'bs-Cyrl', 'bs-Latn', 'de-1901',
	'de-1996', 'de-AT-1901', 'de-AT-1996', 'de-CH-1901', 'de-CH-1996', 'de-DE-1901', 'de-DE-1996',
	'en-boont', 'en-scouse', 'es-419', 'iu-Cans', 'iu-Latn', 'mn-Cyrl', 'mn-Mong', 'sl-nedis',
	'sl-rozaj', 'sr-Cyrl', 'sr-Latn', 'tg-Arab', 'tg-Cyrl', 'uz-Cyrl', 'uz-Latn', 'yi-Latn',
	'zh-Hans', 'zh-Hans-CN', 'zh-Hans-HK', 'zh-Hans-MO', 'zh-Hans-SG', 'zh-Hans-TW', 'zh-Hant',
	'zh-Hant-CN', 'zh-Hant-HK', 'zh-Hant-MO', 'zh-Hant-SG', 'zh-Hant-TW']
