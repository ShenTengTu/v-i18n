module language

pub const variants = ['az-baku1926', 'ba-baku1926', 'be-1959acad', 'be-tarask', 'bg-ivanchov',
	'blo-balanka', 'bo-Latn-pinyin', 'ca-valencia', 'crh-baku1926', 'da-bornholm', 'de-1901',
	'de-1996', 'djk-aluku', 'djk-ndyuka', 'djk-pamaka', 'el-monoton', 'el-polyton', 'en-CA-newfound',
	'en-basiceng', 'en-boont', 'en-cornu', 'en-emodeng', 'en-oxendict', 'en-scotland', 'en-scouse',
	'en-spanglis', 'en-unifon', 'eo-arkaika', 'eo-hsistemo', 'eo-xsistemo', 'es-spanglis',
	'eu-biscayan', 'fr-1694acad', 'frm-1606nict', 'gl-ao1990', 'hnj-pahawh2', 'hnj-pahawh3',
	'hnj-pahawh4', 'hup-unifon', 'ja-Latn-hepburn', 'kea-barla', 'kea-sotav', 'kk-baku1926',
	'kl-tunumiit', 'krc-baku1926', 'kw-kkcor', 'kw-kscor', 'kw-uccor', 'kw-ucrcor', 'ky-baku1926',
	'kyh-unifon', 'la-peano', 'lv-vecdruka', 'mww-pahawh2', 'mww-pahawh3', 'mww-pahawh4',
	'nn-hognorsk', 'oc-aranes', 'oc-aranes-grclass', 'oc-aranes-grmistr', 'oc-auvern',
	'oc-auvern-grclass', 'oc-auvern-grmistr', 'oc-cisaup', 'oc-cisaup-grclass', 'oc-cisaup-grital',
	'oc-cisaup-grmistr', 'oc-creiss', 'oc-creiss-grclass', 'oc-creiss-grmistr', 'oc-gascon',
	'oc-gascon-grclass', 'oc-gascon-grmistr', 'oc-grclass', 'oc-grital', 'oc-grmistr', 'oc-lemosin',
	'oc-lemosin-grclass', 'oc-lemosin-grmistr', 'oc-lengadoc', 'oc-lengadoc-grclass',
	'oc-lengadoc-grmistr', 'oc-nicard', 'oc-nicard-grclass', 'oc-nicard-grital', 'oc-nicard-grmistr',
	'oc-provenc', 'oc-provenc-grclass', 'oc-provenc-grital', 'oc-provenc-grmistr', 'oc-vivaraup',
	'oc-vivaraup-grclass', 'oc-vivaraup-grmistr', 'pl-kociewie', 'pt-BR-abl1943', 'pt-ao1990',
	'pt-colb1945', 'rm-jauer', 'rm-puter', 'rm-rumgr', 'rm-surmiran', 'rm-sursilv', 'rm-sutsilv',
	'rm-vallader', 'ru-luna1918', 'ru-petr1708', 'sa-bauddha', 'sa-itihasa', 'sa-laukika',
	'sa-vaidika', 'sah-baku1926', 'sco-ulster', 'sl-bohoric', 'sl-dajnko', 'sl-metelko', 'sl-nedis',
	'sl-rozaj', 'sl-rozaj-1994', 'sl-rozaj-biske', 'sl-rozaj-biske-1994', 'sl-rozaj-lipaw',
	'sl-rozaj-njiva', 'sl-rozaj-njiva-1994', 'sl-rozaj-osojs', 'sl-rozaj-osojs-1994',
	'sl-rozaj-solba', 'sl-rozaj-solba-1994', 'sr-Cyrl-ekavsk', 'sr-Cyrl-ijekavsk', 'sr-Latn-ekavsk',
	'sr-Latn-ijekavsk', 'sr-ekavsk', 'sr-ijekavsk', 'tk-baku1926', 'tol-unifon', 'tt-baku1926',
	'tw-akuapem', 'tw-asante', 'uz-baku1926', 'vo-nulik', 'vo-rigik', 'yue-jyutping', 'yur-unifon',
	'zh-Latn-pinyin', 'zh-Latn-tongyong', 'zh-Latn-wadegile']
